/*

	Alex Dunker
	adunker@purdue.edu

	Mitch Bouma
	mbouma@purdue.edu

	Hazard Unit

*/

`include "cpu_types_pkg.vh"
`include "hazard_unit_if.vh"

import cpu_types_pkg::*;

module hazard_unit (
	input logic CLK, nRST,
	hazard_unit_if huif
);



endmodule // hazard_unit